module controlUnit(input  logic       clk, reset,
                   input  logic [7:0] instructionByte);



endmodule
