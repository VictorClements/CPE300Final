module smg(input  logic clk, reset, start,
           );
